/****************************************************************************
 *   Copyright (c) 2023 Wenxu Cao
 *  
 *   Filename:         transpose_20.v
 *   Institution:      UESTC
 *   Author:           Wenxu Cao
 *   Version:          1.0
 *   Date:             2023-06-08
 *   Description:      This is a matrix transpose unit.
 *
*****************************************************************************/

module transpose_20(
    input       wire        [19 : 0]        input_0,
    input       wire        [19 : 0]        input_1,
    input       wire        [19 : 0]        input_2,
    input       wire        [19 : 0]        input_3,
    input       wire        [19 : 0]        input_4,
    input       wire        [19 : 0]        input_5,
    input       wire        [19 : 0]        input_6,
    input       wire        [19 : 0]        input_7,
    input       wire        [19 : 0]        input_8,
    input       wire        [19 : 0]        input_9,
    input       wire        [19 : 0]        input_10,
    input       wire        [19 : 0]        input_11,
    input       wire        [19 : 0]        input_12,
    input       wire        [19 : 0]        input_13,
    input       wire        [19 : 0]        input_14,
    input       wire        [19 : 0]        input_15,
    input       wire        [19 : 0]        input_16,
    input       wire        [19 : 0]        input_17,
    input       wire        [19 : 0]        input_18,
    input       wire        [19 : 0]        input_19,

    output      wire        [19 : 0]        output_0,
    output      wire        [19 : 0]        output_1,
    output      wire        [19 : 0]        output_2,
    output      wire        [19 : 0]        output_3,
    output      wire        [19 : 0]        output_4,
    output      wire        [19 : 0]        output_5,
    output      wire        [19 : 0]        output_6,
    output      wire        [19 : 0]        output_7,
    output      wire        [19 : 0]        output_8,
    output      wire        [19 : 0]        output_9,
    output      wire        [19 : 0]        output_10,
    output      wire        [19 : 0]        output_11,
    output      wire        [19 : 0]        output_12,
    output      wire        [19 : 0]        output_13,
    output      wire        [19 : 0]        output_14,
    output      wire        [19 : 0]        output_15,
    output      wire        [19 : 0]        output_16,
    output      wire        [19 : 0]        output_17,
    output      wire        [19 : 0]        output_18,
    output      wire        [19 : 0]        output_19
);

assign output_0 = {
    input_19[0], 
    input_18[0],
    input_17[0],
    input_16[0],
    input_15[0],
    input_14[0],
    input_13[0],
    input_12[0],
    input_11[0],
    input_10[0],
    input_9[0],
    input_8[0],
    input_7[0],
    input_6[0],
    input_5[0],
    input_4[0],
    input_3[0],
    input_2[0],
    input_1[0],
    input_0[0]
};

assign output_1 = {
    input_19[1], 
    input_18[1],
    input_17[1],
    input_16[1],
    input_15[1],
    input_14[1],
    input_13[1],
    input_12[1],
    input_11[1],
    input_10[1],
    input_9[1],
    input_8[1],
    input_7[1],
    input_6[1],
    input_5[1],
    input_4[1],
    input_3[1],
    input_2[1],
    input_1[1],
    input_0[1]
};

assign output_2 = {
    input_19[2], 
    input_18[2],
    input_17[2],
    input_16[2],
    input_15[2],
    input_14[2],
    input_13[2],
    input_12[2],
    input_11[2],
    input_10[2],
    input_9[2],
    input_8[2],
    input_7[2],
    input_6[2],
    input_5[2],
    input_4[2],
    input_3[2],
    input_2[2],
    input_1[2],
    input_0[2]
};

assign output_3 = {
    input_19[3], 
    input_18[3],
    input_17[3],
    input_16[3],
    input_15[3],
    input_14[3],
    input_13[3],
    input_12[3],
    input_11[3],
    input_10[3],
    input_9[3],
    input_8[3],
    input_7[3],
    input_6[3],
    input_5[3],
    input_4[3],
    input_3[3],
    input_2[3],
    input_1[3],
    input_0[3]
};

assign output_4 = {
    input_19[4], 
    input_18[4],
    input_17[4],
    input_16[4],
    input_15[4],
    input_14[4],
    input_13[4],
    input_12[4],
    input_11[4],
    input_10[4],
    input_9[4],
    input_8[4],
    input_7[4],
    input_6[4],
    input_5[4],
    input_4[4],
    input_3[4],
    input_2[4],
    input_1[4],
    input_0[4]
};

assign output_5 = {
    input_19[5], 
    input_18[5],
    input_17[5],
    input_16[5],
    input_15[5],
    input_14[5],
    input_13[5],
    input_12[5],
    input_11[5],
    input_10[5],
    input_9[5],
    input_8[5],
    input_7[5],
    input_6[5],
    input_5[5],
    input_4[5],
    input_3[5],
    input_2[5],
    input_1[5],
    input_0[5]
};

assign output_6 = {
    input_19[6], 
    input_18[6],
    input_17[6],
    input_16[6],
    input_15[6],
    input_14[6],
    input_13[6],
    input_12[6],
    input_11[6],
    input_10[6],
    input_9[6],
    input_8[6],
    input_7[6],
    input_6[6],
    input_5[6],
    input_4[6],
    input_3[6],
    input_2[6],
    input_1[6],
    input_0[6]
};

assign output_7 = {
    input_19[7], 
    input_18[7],
    input_17[7],
    input_16[7],
    input_15[7],
    input_14[7],
    input_13[7],
    input_12[7],
    input_11[7],
    input_10[7],
    input_9[7],
    input_8[7],
    input_7[7],
    input_6[7],
    input_5[7],
    input_4[7],
    input_3[7],
    input_2[7],
    input_1[7],
    input_0[7]
};

assign output_8 = {
    input_19[8], 
    input_18[8],
    input_17[8],
    input_16[8],
    input_15[8],
    input_14[8],
    input_13[8],
    input_12[8],
    input_11[8],
    input_10[8],
    input_9[8],
    input_8[8],
    input_7[8],
    input_6[8],
    input_5[8],
    input_4[8],
    input_3[8],
    input_2[8],
    input_1[8],
    input_0[8]
};

assign output_9 = {
    input_19[9], 
    input_18[9],
    input_17[9],
    input_16[9],
    input_15[9],
    input_14[9],
    input_13[9],
    input_12[9],
    input_11[9],
    input_10[9],
    input_9[9],
    input_8[9],
    input_7[9],
    input_6[9],
    input_5[9],
    input_4[9],
    input_3[9],
    input_2[9],
    input_1[9],
    input_0[9]
};

assign output_10 = {
    input_19[10], 
    input_18[10],
    input_17[10],
    input_16[10],
    input_15[10],
    input_14[10],
    input_13[10],
    input_12[10],
    input_11[10],
    input_10[10],
    input_9[10],
    input_8[10],
    input_7[10],
    input_6[10],
    input_5[10],
    input_4[10],
    input_3[10],
    input_2[10],
    input_1[10],
    input_0[10]
};

assign output_11 = {
    input_19[11], 
    input_18[11],
    input_17[11],
    input_16[11],
    input_15[11],
    input_14[11],
    input_13[11],
    input_12[11],
    input_11[11],
    input_10[11],
    input_9[11],
    input_8[11],
    input_7[11],
    input_6[11],
    input_5[11],
    input_4[11],
    input_3[11],
    input_2[11],
    input_1[11],
    input_0[11]
};

assign output_12 = {
    input_19[12], 
    input_18[12],
    input_17[12],
    input_16[12],
    input_15[12],
    input_14[12],
    input_13[12],
    input_12[12],
    input_11[12],
    input_10[12],
    input_9[12],
    input_8[12],
    input_7[12],
    input_6[12],
    input_5[12],
    input_4[12],
    input_3[12],
    input_2[12],
    input_1[12],
    input_0[12]
};

assign output_13 = {
    input_19[13], 
    input_18[13],
    input_17[13],
    input_16[13],
    input_15[13],
    input_14[13],
    input_13[13],
    input_12[13],
    input_11[13],
    input_10[13],
    input_9[13],
    input_8[13],
    input_7[13],
    input_6[13],
    input_5[13],
    input_4[13],
    input_3[13],
    input_2[13],
    input_1[13],
    input_0[13]
};

assign output_14 = {
    input_19[14], 
    input_18[14],
    input_17[14],
    input_16[14],
    input_15[14],
    input_14[14],
    input_13[14],
    input_12[14],
    input_11[14],
    input_10[14],
    input_9[14],
    input_8[14],
    input_7[14],
    input_6[14],
    input_5[14],
    input_4[14],
    input_3[14],
    input_2[14],
    input_1[14],
    input_0[14]
};

assign output_15 = {
    input_19[15], 
    input_18[15],
    input_17[15],
    input_16[15],
    input_15[15],
    input_14[15],
    input_13[15],
    input_12[15],
    input_11[15],
    input_10[15],
    input_9[15],
    input_8[15],
    input_7[15],
    input_6[15],
    input_5[15],
    input_4[15],
    input_3[15],
    input_2[15],
    input_1[15],
    input_0[15]
};

assign output_16 = {
    input_19[16], 
    input_18[16],
    input_17[16],
    input_16[16],
    input_15[16],
    input_14[16],
    input_13[16],
    input_12[16],
    input_11[16],
    input_10[16],
    input_9[16],
    input_8[16],
    input_7[16],
    input_6[16],
    input_5[16],
    input_4[16],
    input_3[16],
    input_2[16],
    input_1[16],
    input_0[16]
};

assign output_17 = {
    input_19[17], 
    input_18[17],
    input_17[17],
    input_16[17],
    input_15[17],
    input_14[17],
    input_13[17],
    input_12[17],
    input_11[17],
    input_10[17],
    input_9[17],
    input_8[17],
    input_7[17],
    input_6[17],
    input_5[17],
    input_4[17],
    input_3[17],
    input_2[17],
    input_1[17],
    input_0[17]
};

assign output_18 = {
    input_19[18], 
    input_18[18],
    input_17[18],
    input_16[18],
    input_15[18],
    input_14[18],
    input_13[18],
    input_12[18],
    input_11[18],
    input_10[18],
    input_9[18],
    input_8[18],
    input_7[18],
    input_6[18],
    input_5[18],
    input_4[18],
    input_3[18],
    input_2[18],
    input_1[18],
    input_0[18]
};

assign output_19 = {
    input_19[19], 
    input_18[19],
    input_17[19],
    input_16[19],
    input_15[19],
    input_14[19],
    input_13[19],
    input_12[19],
    input_11[19],
    input_10[19],
    input_9[19],
    input_8[19],
    input_7[19],
    input_6[19],
    input_5[19],
    input_4[19],
    input_3[19],
    input_2[19],
    input_1[19],
    input_0[19]
};

endmodule